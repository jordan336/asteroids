library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--Sprite Table
entity sprite_table is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(31 downto 0)
   );
end sprite_table;

architecture arch of sprite_table is
   
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=32;
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
   
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
        
   -- ROM definition
   constant ROM: rom_type:=( 
     -- code x00
   "00000000000000000000000000000000", -- 00
   "00000000000000000000000000000000", -- 01
   "00000000000000000000000000000000", -- 02
   "00000000000000000000000000000000", -- 03
   "00000000000000000000000000000000", -- 04
   "00000000000000000000000000000000", -- 05
   "00000000000000010000000000000000", -- 06                    *
   "00000000000000101000000000000000", -- 07                   * *
   "00000000000001000100000000000000", -- 08                  *   *
   "00000000000010000010000000000000", -- 09                 *     *
   "00000000000100000001000000000000", -- 0a                *       *
   "00000000001000000000100000000000", -- 0b               *         * 
   "00000000010000000000010000000000", -- 0c              *           *
   "00000000100000000000001000000000", -- 0d             *             *
   "00000001000000000000000100000000", -- 0e            *               * 
   "00000010000000000000000010000000", -- 0f           *                 *
   "00000100000000000000000001000000", -- 10          *                   *
   "00001000000000000000000000100000", -- 11         *                     * 
   "00010000000000000000000000010000", -- 12        *                       *
   "00111111111111111111111111111000", -- 13       *************************** 
   "01000000000000000000000000000100", -- 14      *                           * 
   "10000000000000000000000000000010", -- 15     *                             * 
   "00000000000000000000000000000000", -- 16
   "00000000000000000000000000000000", -- 17
   "00000000000000000000000000000000", -- 18
   "00000000000000000000000000000000", -- 19
   "00000000000000000000000000000000", -- 1a
   "00000000000000000000000000000000", -- 1b
   "00000000000000000000000000000000", -- 1c
   "00000000000000000000000000000000", -- 1d
   "00000000000000000000000000000000", -- 1e
   "00000000000000000000000000000000", -- 1f
     -- code x01
   "00000000000000000000000000000000", -- 00
   "00000000000000000000000000000000", -- 01
   "00000000000000000000000000000000", -- 02
   "00000000000000000000000000000000", -- 03
   "00000000000000000000000000000000", -- 04
   "00000000000000000000000000000000", -- 05
   "00000000000000000000000000000000", -- 06
   "00000000000000000000000000000000", -- 07
   "00000000000000000000000000000000", -- 08
   "00000000000000000000000000000000", -- 09
   "00000000000000000000000000000000", -- 0a
   "00000000000000010000000000000000", -- 0b
   "00000000000000111000000000000000", -- 0c
   "00000000000000111000000000000000", -- 0d
   "00000000000000111000000000000000", -- 0e
   "00000000000000010000000000000000", -- 0f
   "00000000000000000000000000000000", -- 10
   "00000000000000000000000000000000", -- 11
   "00000000000000000000000000000000", -- 12
   "00000000000000000000000000000000", -- 13
   "00000000000000000000000000000000", -- 14
   "00000000000000000000000000000000", -- 15
   "00000000000000000000000000000000", -- 16
   "00000000000000000000000000000000", -- 17
   "00000000000000000000000000000000", -- 18
   "00000000000000000000000000000000", -- 19
   "00000000000000000000000000000000", -- 1a
   "00000000000000000000000000000000", -- 1b
   "00000000000000000000000000000000", -- 1c
   "00000000000000000000000000000000", -- 1d
   "00000000000000000000000000000000", -- 1e
   "00000000000000000000000000000000", -- 1f
      -- code x02
   "00000000000000000000000000000000", -- 00
   "00000000000000000000010000000000", -- 01
   "00000000000000000000100000000000", -- 02
   "00000000000000000001000000000000", -- 03
   "00000000000000000011000000000000", -- 04
   "00000000000000000101000000000000", -- 05
   "00000000000000001001000000000000", -- 06
   "00000000000000010001000000000000", -- 07
   "00000000000000100001000000000000", -- 08
   "00000000000001000001000000000000", -- 09
   "00000000000010000001000000000000", -- 0a
   "00000000000100000001000000000000", -- 0b
   "00000000001000000001000000000000", -- 0c
   "00000000010000000001000000000000", -- 0d
   "00000000100000000001000000000000", -- 0e
   "00000001000000000001000000000000", -- 0f
   "00000010000000000001000000000000", -- 10               <
   "00000001000000000001000000000000", -- 11
   "00000000100000000001000000000000", -- 12
   "00000000010000000001000000000000", -- 13
   "00000000001000000001000000000000", -- 14
   "00000000000100000001000000000000", -- 15
   "00000000000010000001000000000000", -- 16
   "00000000000001000001000000000000", -- 17
   "00000000000000100001000000000000", -- 18
   "00000000000000010001000000000000", -- 19
   "00000000000000001001000000000000", -- 1a
   "00000000000000000101000000000000", -- 1b
   "00000000000000000011000000000000", -- 1c
   "00000000000000000001000000000000", -- 1d
   "00000000000000000000100000000000", -- 1e
   "00000000000000000000010000000000", -- 1f
      -- code x03
   "00000000000000000000000000000000", -- 00
   "00000000000000000000000000000000", -- 01
   "00000000000000000000000000000000", -- 02
   "00000000000000000000000000000000", -- 03
   "00000000000000000000000000000000", -- 04
   "00000000000000000000000000000000", -- 05
   "00000000000000000000000000000000", -- 06
   "00000000000000000000000000000000", -- 07
   "00000000000000000000000000000000", -- 08
   "00000000000000000000000000000000", -- 09
   "00000000000000000000000000000000", -- 0a
   "00000000000000010000000000000000", -- 0b
   "00000000000000111000000000000000", -- 0c
   "00000000000000111000000000000000", -- 0d
   "00000000000000111000000000000000", -- 0e
   "00000000000000010000000000000000", -- 0f
   "00000000000000000000000000000000", -- 10
   "00000000000000000000000000000000", -- 11
   "00000000000000000000000000000000", -- 12
   "00000000000000000000000000000000", -- 13
   "00000000000000000000000000000000", -- 14
   "00000000000000000000000000000000", -- 15
   "00000000000000000000000000000000", -- 16
   "00000000000000000000000000000000", -- 17
   "00000000000000000000000000000000", -- 18
   "00000000000000000000000000000000", -- 19
   "00000000000000000000000000000000", -- 1a
   "00000000000000000000000000000000", -- 1b
   "00000000000000000000000000000000", -- 1c
   "00000000000000000000000000000000", -- 1d
   "00000000000000000000000000000000", -- 1e
   "00000000000000000000000000000000", -- 1f
      -- code x04
   "00000000000000000000000000000000", -- 00
   "00000000000000000000000000000000", -- 01
   "00000000000000000000000000000000", -- 02
   "00000000000000000000000000000000", -- 03
   "00000000000000000000000000000000", -- 04
   "00000000000000000000000000000000", -- 05
   "00000000000000000000000000000000", -- 06
   "00000000000000000000000000000000", -- 07
   "00000000000000000000000000000000", -- 08
   "00000000000000000000000000000000", -- 09
   "01000000000000000000000000000001", -- 0a
   "00100000000000000000000000000010", -- 0b
   "00011111111111111111111111111110", -- 0c
   "00001000000000000000000000001000", -- 0d
   "00000100000000000000000000010000", -- 0e
   "00000010000000000000000000100000", -- 0f              \/
   "00000001000000000000000001000000", -- 10
   "00000000100000000000000010000000", -- 11
   "00000000010000000000000100000000", -- 12
   "00000000001000000000001000000000", -- 13
   "00000000000100000000010000000000", -- 14
   "00000000000010000000100000000000", -- 15
   "00000000000001000001000000000000", -- 16
   "00000000000000100010000000000000", -- 17
   "00000000000000010100000000000000", -- 18
   "00000000000000001000000000000000", -- 19
   "00000000000000000000000000000000", -- 1a
   "00000000000000000000000000000000", -- 1b
   "00000000000000000000000000000000", -- 1c
   "00000000000000000000000000000000", -- 1d
   "00000000000000000000000000000000", -- 1e
   "00000000000000000000000000000000", -- 1f
      -- code x05
   "00000000000000000000000000000000", -- 00
   "00000000000000000000000000000000", -- 01
   "00000000000000000000000000000000", -- 02
   "00000000000000000000000000000000", -- 03
   "00000000000000000000000000000000", -- 04
   "00000000000000000000000000000000", -- 05
   "00000000000000000000000000000000", -- 06
   "00000000000000000000000000000000", -- 07
   "00000000000000000000000000000000", -- 08
   "00000000000000000000000000000000", -- 09
   "00000000000000000000000000000000", -- 0a
   "00000000000000010000000000000000", -- 0b
   "00000000000000111000000000000000", -- 0c
   "00000000000000111000000000000000", -- 0d
   "00000000000000111000000000000000", -- 0e
   "00000000000000010000000000000000", -- 0f
   "00000000000000000000000000000000", -- 10
   "00000000000000000000000000000000", -- 11
   "00000000000000000000000000000000", -- 12
   "00000000000000000000000000000000", -- 13
   "00000000000000000000000000000000", -- 14
   "00000000000000000000000000000000", -- 15
   "00000000000000000000000000000000", -- 16
   "00000000000000000000000000000000", -- 17
   "00000000000000000000000000000000", -- 18
   "00000000000000000000000000000000", -- 19
   "00000000000000000000000000000000", -- 1a
   "00000000000000000000000000000000", -- 1b
   "00000000000000000000000000000000", -- 1c
   "00000000000000000000000000000000", -- 1d
   "00000000000000000000000000000000", -- 1e
   "00000000000000000000000000000000", -- 1f
      -- code x06
   "00000000001000000000000000000000", -- 00
   "00000000000100000000000000000000", -- 01
   "00000000000010000000000000000000", -- 02
   "00000000000011000000000000000000", -- 03
   "00000000000010100000000000000000", -- 04
   "00000000000010010000000000000000", -- 05
   "00000000000010001000000000000000", -- 06
   "00000000000010000100000000000000", -- 07
   "00000000000010000010000000000000", -- 08
   "00000000000010000001000000000000", -- 09
   "00000000000010000000100000000000", -- 0a
   "00000000000010000000010000000000", -- 0b
   "00000000000010000000001000000000", -- 0c
   "00000000000010000000000100000000", -- 0d
   "00000000000010000000000010000000", -- 0e              >
   "00000000000010000000000001000000", -- 0f
   "00000000000010000000000010000000", -- 10
   "00000000000010000000000100000000", -- 11
   "00000000000010000000001000000000", -- 12
   "00000000000010000000010000000000", -- 13
   "00000000000010000000100000000000", -- 14
   "00000000000010000001000000000000", -- 15
   "00000000000010000010000000000000", -- 16
   "00000000000010000100000000000000", -- 17
   "00000000000010001000000000000000", -- 18
   "00000000000010010000000000000000", -- 19
   "00000000000010100000000000000000", -- 1a
   "00000000000011000000000000000000", -- 1b
   "00000000000010000000000000000000", -- 1c
   "00000000000100000000000000000000", -- 1d
   "00000000001000000000000000000000", -- 1e
   "00000000000000000000000000000000", -- 1f
         -- code x07
   "00000000000000000000000000000000", -- 00
   "00000000000000000000000000000000", -- 01
   "00000000000000000000000000000000", -- 02
   "00000000000000000000000000000000", -- 03
   "00000000000000000000000000000000", -- 04
   "00000000000000000000000000000000", -- 05
   "00000000000000000000000000000000", -- 06
   "00000000000000000000000000000000", -- 07
   "00000000000000000000000000000000", -- 08
   "00000000000000000000000000000000", -- 09
   "00000000000000000000000000000000", -- 0a
   "00000000000000000000000000000000", -- 0b
   "00000000000000011100000000000000", -- 0c
   "00000000000000011100000000000000", -- 0d
   "00000000000011111111100000000000", -- 0e
   "00000000000011111111100000000000", -- 0f
   "00000000000000011100000000000000", -- 10
   "00000000000000011100000000000000", -- 11
   "00000000000000000000000000000000", -- 12
   "00000000000000000000000000000000", -- 13
   "00000000000000000000000000000000", -- 14
   "00000000000000000000000000000000", -- 15
   "00000000000000000000000000000000", -- 16
   "00000000000000000000000000000000", -- 17
   "00000000000000000000000000000000", -- 18
   "00000000000000000000000000000000", -- 19
   "00000000000000000000000000000000", -- 1a
   "00000000000000000000000000000000", -- 1b
   "00000000000000000000000000000000", -- 1c
   "00000000000000000000000000000000", -- 1d
   "00000000000000000000000000000000", -- 1e
   "00000000000000000000000000000000"  -- 1f
   );
      
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        addr_reg <= addr;
      end if;
   end process;
   data <= ROM(to_integer(unsigned(addr_reg)));
end arch;
